Amplitudovy modulator s AD633
*
.LIB AD633.lib
*
.PARAM nosna_f=50k
.PARAM modulovana_f=1k
*
XAM X1 0 Y1 0 VNEG Y1 W VPOS ad633; AD633
* modulovaný a nosný vstupný signál
Vm X1 0 AC 1 0 SIN(0 1 {modulovana_f})
Vn Y1 0 AC 15 0 SIN(0 1 {nosna_f})
* napájanie
Vpos VPOS 0 15V
Vneg VNEG 0 -15V

C1 VPOS 0 0.1u
C2 VNEG 0 0.1u
*
.TRAN 1u 1m
.PROBE V(W,0) V(X1,0) V(Y1,0)

.END
